# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xnor2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 5.930000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.075000 2.005000 1.275000 ;
        RECT 1.835000 1.275000 2.005000 1.445000 ;
        RECT 1.835000 1.445000 6.270000 1.615000 ;
        RECT 6.100000 1.075000 8.170000 1.275000 ;
        RECT 6.100000 1.275000 6.270000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.858500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  6.750000 1.785000  9.060000 2.045000 ;
        RECT  8.730000 1.445000 10.940000 1.665000 ;
        RECT  8.730000 1.665000  9.060000 1.785000 ;
        RECT  8.730000 2.045000  9.060000 2.465000 ;
        RECT  9.150000 0.655000 10.940000 0.905000 ;
        RECT  9.710000 1.665000  9.960000 2.465000 ;
        RECT 10.610000 1.665000 10.940000 2.465000 ;
        RECT 10.705000 0.905000 10.940000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.645000  1.910000 0.905000 ;
      RECT  0.085000  0.905000  0.320000 1.445000 ;
      RECT  0.085000  1.445000  1.400000 1.615000 ;
      RECT  0.085000  1.615000  0.460000 2.465000 ;
      RECT  0.170000  0.255000  2.380000 0.475000 ;
      RECT  0.680000  1.835000  0.930000 2.635000 ;
      RECT  1.150000  1.615000  1.400000 1.785000 ;
      RECT  1.150000  1.785000  4.220000 2.005000 ;
      RECT  1.150000  2.005000  1.400000 2.465000 ;
      RECT  1.620000  2.175000  1.870000 2.635000 ;
      RECT  2.090000  2.005000  2.340000 2.465000 ;
      RECT  2.130000  0.475000  2.380000 0.725000 ;
      RECT  2.130000  0.725000  4.260000 0.905000 ;
      RECT  2.560000  2.175000  2.810000 2.635000 ;
      RECT  2.600000  0.085000  2.770000 0.555000 ;
      RECT  2.940000  0.255000  3.320000 0.725000 ;
      RECT  3.030000  2.005000  3.280000 2.465000 ;
      RECT  3.500000  2.175000  3.750000 2.635000 ;
      RECT  3.540000  0.085000  3.710000 0.555000 ;
      RECT  3.880000  0.255000  4.260000 0.725000 ;
      RECT  3.970000  2.005000  4.220000 2.465000 ;
      RECT  4.425000  1.785000  6.580000 2.005000 ;
      RECT  4.425000  2.005000  4.740000 2.465000 ;
      RECT  4.430000  0.085000  4.700000 0.905000 ;
      RECT  4.870000  0.255000  5.250000 0.725000 ;
      RECT  4.870000  0.725000  8.170000 0.735000 ;
      RECT  4.870000  0.735000  8.980000 0.905000 ;
      RECT  4.960000  2.175000  5.210000 2.635000 ;
      RECT  5.430000  2.005000  5.680000 2.465000 ;
      RECT  5.470000  0.085000  5.640000 0.555000 ;
      RECT  5.810000  0.255000  6.190000 0.725000 ;
      RECT  5.900000  2.175000  6.150000 2.635000 ;
      RECT  6.370000  2.005000  6.580000 2.215000 ;
      RECT  6.370000  2.215000  8.540000 2.465000 ;
      RECT  6.410000  0.085000  6.580000 0.555000 ;
      RECT  6.490000  1.445000  8.560000 1.615000 ;
      RECT  6.750000  0.255000  7.130000 0.725000 ;
      RECT  7.350000  0.085000  7.520000 0.555000 ;
      RECT  7.690000  0.255000  8.070000 0.725000 ;
      RECT  8.290000  0.085000  8.460000 0.555000 ;
      RECT  8.390000  1.075000 10.535000 1.275000 ;
      RECT  8.390000  1.275000  8.560000 1.445000 ;
      RECT  8.730000  0.305000 10.940000 0.475000 ;
      RECT  8.730000  0.475000  8.980000 0.735000 ;
      RECT  9.240000  1.835000  9.490000 2.635000 ;
      RECT 10.180000  1.835000 10.430000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.165000  1.445000  1.335000 1.615000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.725000  1.445000  6.895000 1.615000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 1.055000 1.415000 1.395000 1.460000 ;
      RECT 1.055000 1.460000 7.005000 1.600000 ;
      RECT 1.055000 1.600000 1.395000 1.645000 ;
      RECT 6.655000 1.415000 7.005000 1.460000 ;
      RECT 6.655000 1.600000 7.005000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_4
END LIBRARY
