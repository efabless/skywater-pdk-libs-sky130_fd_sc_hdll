# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__bufinv_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.505000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 0.260000 3.295000 0.735000 ;
        RECT 2.915000 0.735000 6.805000 0.905000 ;
        RECT 2.915000 1.445000 6.805000 1.615000 ;
        RECT 2.915000 1.615000 3.295000 2.465000 ;
        RECT 3.855000 0.260000 4.235000 0.735000 ;
        RECT 3.855000 1.615000 4.235000 2.465000 ;
        RECT 4.795000 0.260000 5.175000 0.735000 ;
        RECT 4.795000 1.615000 5.175000 2.465000 ;
        RECT 5.735000 0.260000 6.115000 0.735000 ;
        RECT 5.735000 1.615000 6.115000 2.465000 ;
        RECT 6.415000 0.905000 6.805000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.260000 0.895000 0.905000 ;
      RECT 0.515000  1.545000 0.895000 2.465000 ;
      RECT 0.725000  0.905000 0.895000 1.075000 ;
      RECT 0.725000  1.075000 2.355000 1.275000 ;
      RECT 0.725000  1.275000 0.895000 1.545000 ;
      RECT 1.085000  0.260000 1.415000 0.735000 ;
      RECT 1.085000  0.735000 2.745000 0.905000 ;
      RECT 1.085000  1.445000 2.745000 1.615000 ;
      RECT 1.085000  1.615000 1.415000 2.465000 ;
      RECT 1.635000  0.085000 1.805000 0.565000 ;
      RECT 1.635000  1.785000 1.805000 2.635000 ;
      RECT 1.975000  0.260000 2.355000 0.735000 ;
      RECT 1.975000  1.615000 2.355000 2.465000 ;
      RECT 2.575000  0.085000 2.745000 0.565000 ;
      RECT 2.575000  0.905000 2.745000 1.075000 ;
      RECT 2.575000  1.075000 6.245000 1.275000 ;
      RECT 2.575000  1.275000 2.745000 1.445000 ;
      RECT 2.575000  1.785000 2.745000 2.635000 ;
      RECT 3.515000  0.085000 3.685000 0.565000 ;
      RECT 3.515000  1.835000 3.685000 2.635000 ;
      RECT 4.455000  0.085000 4.625000 0.565000 ;
      RECT 4.455000  1.835000 4.625000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.565000 ;
      RECT 5.395000  1.835000 5.565000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.565000 ;
      RECT 6.335000  1.835000 6.505000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufinv_8
END LIBRARY
