# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  16.10000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.405000 1.075000 3.795000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.245000 1.075000 7.635000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.445000 1.075000 11.835000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.985000 1.075000 15.355000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 0.255000  0.895000 0.725000 ;
        RECT  0.565000 0.725000 15.515000 0.905000 ;
        RECT  1.505000 0.255000  1.835000 0.725000 ;
        RECT  2.445000 0.255000  2.775000 0.725000 ;
        RECT  3.385000 0.255000  3.715000 0.725000 ;
        RECT  4.325000 0.255000  4.655000 0.725000 ;
        RECT  5.265000 0.255000  5.595000 0.725000 ;
        RECT  6.205000 0.255000  6.535000 0.725000 ;
        RECT  7.145000 0.255000  7.475000 0.725000 ;
        RECT  8.605000 0.255000  8.935000 0.725000 ;
        RECT  9.545000 0.255000  9.875000 0.725000 ;
        RECT 10.485000 0.255000 10.815000 0.725000 ;
        RECT 11.425000 0.255000 11.755000 0.725000 ;
        RECT 12.365000 0.255000 12.695000 0.725000 ;
        RECT 12.405000 0.905000 12.815000 1.455000 ;
        RECT 12.405000 1.455000 15.475000 1.625000 ;
        RECT 12.405000 1.625000 12.655000 2.125000 ;
        RECT 13.305000 0.255000 13.635000 0.725000 ;
        RECT 13.345000 1.625000 13.595000 2.125000 ;
        RECT 14.245000 0.255000 14.575000 0.725000 ;
        RECT 14.285000 1.625000 14.535000 2.125000 ;
        RECT 15.185000 0.255000 15.515000 0.725000 ;
        RECT 15.225000 1.625000 15.475000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.100000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.100000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.100000 0.085000 ;
      RECT  0.000000  2.635000 16.100000 2.805000 ;
      RECT  0.095000  1.455000  4.145000 1.625000 ;
      RECT  0.095000  1.625000  0.425000 2.465000 ;
      RECT  0.135000  0.085000  0.395000 0.905000 ;
      RECT  0.605000  1.795000  0.855000 2.635000 ;
      RECT  1.065000  0.085000  1.335000 0.555000 ;
      RECT  1.075000  1.625000  1.325000 2.465000 ;
      RECT  1.545000  1.795000  1.795000 2.635000 ;
      RECT  2.005000  0.085000  2.275000 0.555000 ;
      RECT  2.015000  1.625000  2.265000 2.465000 ;
      RECT  2.485000  1.795000  2.735000 2.635000 ;
      RECT  2.945000  0.085000  3.215000 0.555000 ;
      RECT  2.955000  1.625000  3.205000 2.465000 ;
      RECT  3.425000  1.795000  3.675000 2.635000 ;
      RECT  3.885000  0.085000  4.155000 0.555000 ;
      RECT  3.895000  1.625000  4.145000 2.295000 ;
      RECT  3.895000  2.295000  7.945000 2.465000 ;
      RECT  4.365000  1.455000 11.715000 1.625000 ;
      RECT  4.365000  1.625000  4.615000 2.125000 ;
      RECT  4.825000  0.085000  5.095000 0.555000 ;
      RECT  4.835000  1.795000  5.085000 2.295000 ;
      RECT  5.305000  1.625000  5.555000 2.125000 ;
      RECT  5.765000  0.085000  6.035000 0.555000 ;
      RECT  5.775000  1.795000  6.025000 2.295000 ;
      RECT  6.245000  1.625000  6.495000 2.125000 ;
      RECT  6.705000  0.085000  6.975000 0.555000 ;
      RECT  6.715000  1.795000  6.965000 2.295000 ;
      RECT  7.185000  1.625000  7.435000 2.125000 ;
      RECT  7.645000  0.085000  8.435000 0.555000 ;
      RECT  7.655000  1.795000  7.945000 2.295000 ;
      RECT  8.135000  1.795000  8.425000 2.295000 ;
      RECT  8.135000  2.295000 15.995000 2.465000 ;
      RECT  8.645000  1.625000  8.895000 2.125000 ;
      RECT  9.075000  1.795000  9.365000 2.295000 ;
      RECT  9.105000  0.085000  9.375000 0.555000 ;
      RECT  9.585000  1.625000  9.835000 2.125000 ;
      RECT 10.045000  0.085000 10.315000 0.555000 ;
      RECT 10.055000  1.795000 10.305000 2.295000 ;
      RECT 10.525000  1.625000 10.775000 2.125000 ;
      RECT 10.985000  0.085000 11.255000 0.555000 ;
      RECT 10.995000  1.795000 11.245000 2.295000 ;
      RECT 11.465000  1.625000 11.715000 2.125000 ;
      RECT 11.925000  0.085000 12.195000 0.555000 ;
      RECT 11.935000  1.455000 12.185000 2.295000 ;
      RECT 12.865000  0.085000 13.135000 0.555000 ;
      RECT 12.875000  1.795000 13.125000 2.295000 ;
      RECT 13.805000  0.085000 14.075000 0.555000 ;
      RECT 13.815000  1.795000 14.065000 2.295000 ;
      RECT 14.745000  0.085000 15.015000 0.555000 ;
      RECT 14.755000  1.795000 15.005000 2.295000 ;
      RECT 15.685000  0.085000 15.965000 0.905000 ;
      RECT 15.695000  1.465000 15.995000 2.295000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_8
END LIBRARY
