# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand4b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.180000 1.075000 5.040000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.240000 1.075000 7.110000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.665000 1.075000 9.505000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.736000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 2.840000 0.905000 ;
        RECT 1.505000 1.445000 8.985000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.410000 0.905000 2.840000 1.445000 ;
        RECT 2.445000 1.665000 2.825000 2.465000 ;
        RECT 3.385000 1.665000 3.765000 2.465000 ;
        RECT 4.325000 1.665000 4.705000 2.465000 ;
        RECT 5.785000 1.665000 6.165000 2.465000 ;
        RECT 6.725000 1.665000 7.105000 2.465000 ;
        RECT 7.665000 1.665000 8.045000 2.465000 ;
        RECT 8.605000 1.665000 8.985000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 0.855000 0.905000 ;
      RECT 0.090000  1.495000 0.855000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.895000 0.545000 ;
      RECT 0.645000  1.835000 1.335000 2.635000 ;
      RECT 0.660000  0.905000 0.855000 1.075000 ;
      RECT 0.660000  1.075000 1.975000 1.275000 ;
      RECT 0.660000  1.275000 0.855000 1.495000 ;
      RECT 1.045000  1.495000 1.335000 1.835000 ;
      RECT 1.085000  0.255000 5.175000 0.465000 ;
      RECT 1.085000  0.465000 1.335000 0.905000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 3.045000  1.835000 3.215000 2.635000 ;
      RECT 3.385000  0.635000 7.105000 0.905000 ;
      RECT 3.985000  1.835000 4.155000 2.635000 ;
      RECT 4.925000  1.835000 5.615000 2.635000 ;
      RECT 5.365000  0.255000 7.575000 0.465000 ;
      RECT 6.385000  1.835000 6.555000 2.635000 ;
      RECT 7.325000  0.465000 7.575000 0.735000 ;
      RECT 7.325000  0.735000 9.460000 0.905000 ;
      RECT 7.325000  1.835000 7.495000 2.635000 ;
      RECT 7.795000  0.085000 7.965000 0.545000 ;
      RECT 8.135000  0.255000 8.515000 0.735000 ;
      RECT 8.265000  1.835000 8.435000 2.635000 ;
      RECT 8.735000  0.085000 8.905000 0.545000 ;
      RECT 9.075000  0.255000 9.460000 0.735000 ;
      RECT 9.205000  1.445000 9.460000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_4
END LIBRARY
