* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*
* Updated May 2, 2024 with subcircuit compatible with continuous models

.subckt sky130_fd_sc_hdll__diode_4 DIODE VGND VNB VPB VPWR
XD0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=9.88e+06 area=1.0557e+12
.ends
