/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HDLL__MUXB4TO1_4_PP_BLACKBOX_V
`define SKY130_FD_SC_HDLL__MUXB4TO1_4_PP_BLACKBOX_V

/**
 * muxb4to1: Buffered 4-input multiplexer.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_sc_hdll__muxb4to1_4 (
    Z   ,
    D   ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output       Z   ;
    input  [3:0] D   ;
    input  [3:0] S   ;
    input        VPWR;
    input        VGND;
    input        VPB ;
    input        VNB ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HDLL__MUXB4TO1_4_PP_BLACKBOX_V
